-- ===================================================================================================================================
-- @ Author: Krzysztof Pierczyk
-- @ Create Time: 2021-05-24 02:18:50
-- @ Modified time: 2021-05-24 02:20:16
-- @ Description: 
--    
--    Common generator's package
--    
-- ===================================================================================================================================


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package generator is

    -- Quadruplet generator's mode
    type SIGNESS is (SIGNED_OUT, UNSIGNED_OUT);

end package generator;
