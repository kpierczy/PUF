��- -   T h i s   i s   P a c k a g e   S T A N D A R D   a s   d e f i n e d   i n   t h e   V H D L   2 0 0 8   L a n g u a g e   R e f e r e n c e   M a n u a l .  
 - -  
 - -       N O T E :   V C O M   a n d   V S I M   w i l l   n o t   w o r k   p r o p e r l y   i f   t h e s e   d e c l a r a t i o n s  
 - -                   a r e   m o d i f i e d .  
  
 - -   V e r s i o n   i n f o r m a t i o n :    
 ( # ) s t a n d a r d . v h d 	  
  
 p a c k a g e   S T A N D A R D   i s    
 	 t y p e   B O O L E A N   i s   ( F A L S E , T R U E ) ;    
 	 t y p e   B I T   i s   ( ' 0 ' ,   ' 1 ' ) ;    
 	 t y p e   C H A R A C T E R   i s   (  
 	 	 N U L ,   S O H ,   S T X ,   E T X ,   E O T ,   E N Q ,   A C K ,   B E L ,    
 	 	 B S ,     H T ,     L F ,     V T ,     F F ,     C R ,     S O ,     S I ,    
 	 	 D L E ,   D C 1 ,   D C 2 ,   D C 3 ,   D C 4 ,   N A K ,   S Y N ,   E T B ,    
 	 	 C A N ,   E M ,     S U B ,   E S C ,   F S P ,   G S P ,   R S P ,   U S P ,    
  
 	 	 '   ' ,   ' ! ' ,   ' " ' ,   ' # ' ,   ' $ ' ,   ' % ' ,   ' & ' ,   ' ' ' ,    
 	 	 ' ( ' ,   ' ) ' ,   ' * ' ,   ' + ' ,   ' , ' ,   ' - ' ,   ' . ' ,   ' / ' ,    
 	 	 ' 0 ' ,   ' 1 ' ,   ' 2 ' ,   ' 3 ' ,   ' 4 ' ,   ' 5 ' ,   ' 6 ' ,   ' 7 ' ,    
 	 	 ' 8 ' ,   ' 9 ' ,   ' : ' ,   ' ; ' ,   ' < ' ,   ' = ' ,   ' > ' ,   ' ? ' ,    
  
 	 	 ' @ ' ,   ' A ' ,   ' B ' ,   ' C ' ,   ' D ' ,   ' E ' ,   ' F ' ,   ' G ' ,    
 	 	 ' H ' ,   ' I ' ,   ' J ' ,   ' K ' ,   ' L ' ,   ' M ' ,   ' N ' ,   ' O ' ,    
 	 	 ' P ' ,   ' Q ' ,   ' R ' ,   ' S ' ,   ' T ' ,   ' U ' ,   ' V ' ,   ' W ' ,    
 	 	 ' X ' ,   ' Y ' ,   ' Z ' ,   ' [ ' ,   ' \ ' ,   ' ] ' ,   ' ^ ' ,   ' _ ' ,    
  
 	 	 ' ` ' ,   ' a ' ,   ' b ' ,   ' c ' ,   ' d ' ,   ' e ' ,   ' f ' ,   ' g ' ,    
 	 	 ' h ' ,   ' i ' ,   ' j ' ,   ' k ' ,   ' l ' ,   ' m ' ,   ' n ' ,   ' o ' ,    
 	 	 ' p ' ,   ' q ' ,   ' r ' ,   ' s ' ,   ' t ' ,   ' u ' ,   ' v ' ,   ' w ' ,    
 	 	 ' x ' ,   ' y ' ,   ' z ' ,   ' { ' ,   ' | ' ,   ' } ' ,   ' ~ ' ,   D E L ,  
  
 	 	 C 1 2 8 ,   C 1 2 9 ,   C 1 3 0 ,   C 1 3 1 ,   C 1 3 2 ,   C 1 3 3 ,   C 1 3 4 ,   C 1 3 5 ,  
 	 	 C 1 3 6 ,   C 1 3 7 ,   C 1 3 8 ,   C 1 3 9 ,   C 1 4 0 ,   C 1 4 1 ,   C 1 4 2 ,   C 1 4 3 ,  
 	 	 C 1 4 4 ,   C 1 4 5 ,   C 1 4 6 ,   C 1 4 7 ,   C 1 4 8 ,   C 1 4 9 ,   C 1 5 0 ,   C 1 5 1 ,  
 	 	 C 1 5 2 ,   C 1 5 3 ,   C 1 5 4 ,   C 1 5 5 ,   C 1 5 6 ,   C 1 5 7 ,   C 1 5 8 ,   C 1 5 9 ,  
  
 	 	 - -   t h e   c h a r a c t e r   c o d e   f o r   1 6 0   i s   t h e r e   ( N B S P ) ,    
 	 	 - -   b u t   p r i n t s   a s   n o   c h a r    
  
 	 	 ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,  
 	 	 ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,  
 	 	 ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,  
 	 	 ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,  
  
 	 	 ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,  
 	 	 ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,  
 	 	 ' � ' ,   ' � ' ,   ' � ' ,   ' o ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,  
 	 	 ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,  
  
 	 	 ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,  
 	 	 ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,  
 	 	 ' � ' ,   ' � ' ,   ' � ' ,   ' o ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,  
 	 	 ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � ' ,   ' � '   ) ;    
  
 	 t y p e   S E V E R I T Y _ L E V E L   i s   ( N O T E ,   W A R N I N G ,   E R R O R ,   F A I L U R E ) ;    
 	 t y p e   I N T E G E R   i s   r a n g e   - 2 1 4 7 4 8 3 6 4 8   t o   2 1 4 7 4 8 3 6 4 7 ;    
 	 t y p e   R E A L   i s   r a n g e   - 1 . 0 E 3 0 8   t o   1 . 0 E 3 0 8 ;    
 	 t y p e   T I M E   i s   r a n g e   - 2 1 4 7 4 8 3 6 4 7   t o   2 1 4 7 4 8 3 6 4 7    
 	 	 u n i t s    
 	 	 	 f s ;  
 	 	 	 p s   =   1 0 0 0   f s ;  
 	 	 	 n s   =   1 0 0 0   p s ;  
 	 	 	 u s   =   1 0 0 0   n s ;    
 	 	 	 m s   =   1 0 0 0   u s ;    
 	 	 	 s e c   =   1 0 0 0   m s ;    
 	 	 	 m i n   =   6 0   s e c ;    
 	 	 	 h r   =   6 0   m i n ;    
 	 	 e n d   u n i t s ;  
 	 t y p e   d o m a i n _ t y p e   i s   ( q u i e s c e n t _ d o m a i n ,   t i m e _ d o m a i n ,   f r e q u e n c y _ d o m a i n ) ;   - -   T O D O _ A M S :   A d d   p r e d e f i n e d   o p e r a t o r s  
 	 s i g n a l   d o m a i n :   d o m a i n _ t y p e : = q u i e s c e n t _ d o m a i n ;  
 	 s u b t y p e   D E L A Y _ L E N G T H   i s   T I M E   r a n g e   0   f s   t o   T I M E ' H I G H ;  
 	 i m p u r e   f u n c t i o n   N O W   r e t u r n   D E L A Y _ L E N G T H ;    
 	 i m p u r e   f u n c t i o n   n o w   r e t u r n   r e a l ;  
 	 - -   T O D O _ A M S   - -   f u n c t i o n   f r e q u e n c y   r e t u r n   r e a l ;  
 	 s u b t y p e   N A T U R A L   i s   I N T E G E R   r a n g e   0   t o   I N T E G E R ' H I G H ;    
 	 s u b t y p e   P O S I T I V E   i s   I N T E G E R   r a n g e   1   t o   I N T E G E R ' H I G H ;    
 	 t y p e   S T R I N G   i s   a r r a y   ( P O S I T I V E   r a n g e   < > )   o f   C H A R A C T E R ;    
 	 t y p e   B O O L E A N _ V E C T O R   i s   a r r a y   ( N A T U R A L   r a n g e   < > )   o f   B O O L E A N ;    
 	 t y p e   B I T _ V E C T O R   i s   a r r a y   ( N A T U R A L   r a n g e   < > )   o f   B I T ;    
 	 t y p e   I N T E G E R _ V E C T O R   i s   a r r a y   ( N A T U R A L   r a n g e   < > )   o f   I N T E G E R ;    
 	 t y p e   R E A L _ V E C T O R   i s   a r r a y   ( N A T U R A L   r a n g e   < > )   o f   R E A L ;    
 	 t y p e   T I M E _ V E C T O R   i s   a r r a y   ( N A T U R A L   r a n g e   < > )   o f   T I M E ;    
 	 t y p e   F I L E _ O P E N _ K I N D   i s   (  
 	 	 R E A D _ M O D E ,  
 	 	 W R I T E _ M O D E ,  
 	 	 A P P E N D _ M O D E ) ;  
 	 t y p e   F I L E _ O P E N _ S T A T U S   i s   (  
 	 	 O P E N _ O K ,  
 	 	 S T A T U S _ E R R O R ,  
 	 	 N A M E _ E R R O R ,  
 	 	 M O D E _ E R R O R ) ;  
 	 a t t r i b u t e   F O R E I G N   :   S T R I N G ;  
 e n d   S T A N D A R D ;   