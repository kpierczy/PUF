-- ===================================================================================================================================
-- @ Author: Krzysztof Pierczyk
-- @ Create Time: 2021-04-26 18:18:27
-- @ Modified time: 2021-04-26 18:20:05
-- @ Description:
-- 
--     Uart receiver package's testbench 
--
-- ===================================================================================================================================

library ieee;
use ieee.std_logic_1164.all;
library work;
use work.uart.all;
use work.sim.all;

-- ------------------------------------------------------------- Entity --------------------------------------------------------------

entity uart_rx_tb is
end entity uart_rx_tb;

-- ---------------------------------------------------------- Architecture -----------------------------------------------------------

architecture logic of uart_rx_tb is  
begin
    
    process is
    begin
        wait for 10ns;
    end process;
    
end architecture logic;
